import "DPI-C"
function void bluenoc_recv_tcp_beat( output bit[135:0] result_value
			       , input int unsigned  socket_descriptor
			       , byte         beat_size
			       , byte         bytes_already_received
			       , bit[127:0]   beat_value_so_far
			       );

import "DPI-C"
function byte bluenoc_send_tcp_beat( int unsigned  socket_descriptor
				    , byte          beat_size
				    , byte          bytes_to_send
				    , bit[127:0]    beat_value
				    );

import "DPI-C"
function int unsigned bluenoc_open_tcp_socket( int unsigned tcp_port );
//
// Generated by Bluespec Compiler, version 2017.07.A (build e1df8052c, 2017-07-21)
//
//
//
//
// Ports:
// Name                         I/O  size props
// axi_in_tready                  O     1
// CLK_aclk                       I     1 clock
// RST_N_aresetn                  I     1 reset
// axi_in_tvalid                  I     1
// axi_in_tdata                   I   608 reg
// axi_in_tstrb                   I    76 reg
// axi_in_tkeep                   I    76 reg
// axi_in_tlast                   I     1 reg
// tvswitch                       I     2 reg
//
// No combinational paths from inputs to outputs
//
//

`ifdef BSV_ASSIGNMENT_DELAY
`else
  `define BSV_ASSIGNMENT_DELAY
`endif

`ifdef BSV_POSITIVE_RESET
  `define BSV_RESET_VALUE 1'b1
  `define BSV_RESET_EDGE posedge
`else
  `define BSV_RESET_VALUE 1'b0
  `define BSV_RESET_EDGE negedge
`endif

module mkSVF_Bridge(CLK_aclk,
		    RST_N_aresetn,

		    axi_in_tvalid,
		    axi_in_tdata,
		    axi_in_tstrb,
		    axi_in_tkeep,
		    axi_in_tlast,

		    axi_in_tready,

		    tvswitch);
  input  CLK_aclk;
  input  RST_N_aresetn;

  // action method axi_in_m_tvalid
  input  axi_in_tvalid;
  input  [607 : 0] axi_in_tdata;
  input  [75 : 0] axi_in_tstrb;
  input  [75 : 0] axi_in_tkeep;
  input  axi_in_tlast;

  // value method axi_in_m_tready
  output axi_in_tready;

  // action method tv_switch
  input  [1 : 0] tvswitch;

  // signals for module outputs
  wire axi_in_tready;

  // inlined wires
  wire fOut_dst_ok$wget;

  // register bridge_inReset_isInReset
  reg bridge_inReset_isInReset;
  wire bridge_inReset_isInReset$D_IN, bridge_inReset_isInReset$EN;

  // register bridge_rBeatFromTCP
  reg [31 : 0] bridge_rBeatFromTCP;
  wire [31 : 0] bridge_rBeatFromTCP$D_IN;
  wire bridge_rBeatFromTCP$EN;

  // register bridge_rBeatToTCP
  reg [31 : 0] bridge_rBeatToTCP;
  wire [31 : 0] bridge_rBeatToTCP$D_IN;
  wire bridge_rBeatToTCP$EN;

  // register bridge_rBytesFromTCP
  reg [7 : 0] bridge_rBytesFromTCP;
  wire [7 : 0] bridge_rBytesFromTCP$D_IN;
  wire bridge_rBytesFromTCP$EN;

  // register bridge_rBytesToTCP
  reg [7 : 0] bridge_rBytesToTCP;
  wire [7 : 0] bridge_rBytesToTCP$D_IN;
  wire bridge_rBytesToTCP$EN;

  // register bridge_rFileHandle
  reg [31 : 0] bridge_rFileHandle;
  wire [31 : 0] bridge_rFileHandle$D_IN;
  wire bridge_rFileHandle$EN;

  // register cnt
  reg [7 : 0] cnt;
  wire [7 : 0] cnt$D_IN;
  wire cnt$EN;

  // register trace
  reg [575 : 0] trace;
  wire [575 : 0] trace$D_IN;
  wire trace$EN;

  // register tracesOn
  reg tracesOn;
  wire tracesOn$D_IN, tracesOn$EN;

  // register vecSize
  reg [7 : 0] vecSize;
  wire [7 : 0] vecSize$D_IN;
  wire vecSize$EN;

  // register vrgs_0
  reg [1 : 0] vrgs_0;
  wire [1 : 0] vrgs_0$D_IN;
  wire vrgs_0$EN;

  // register vrgs_1
  reg [1 : 0] vrgs_1;
  wire [1 : 0] vrgs_1$D_IN;
  wire vrgs_1$EN;

  // register vrgs_2
  reg [1 : 0] vrgs_2;
  wire [1 : 0] vrgs_2$D_IN;
  wire vrgs_2$EN;

  // register vrgs_3
  reg [1 : 0] vrgs_3;
  wire [1 : 0] vrgs_3$D_IN;
  wire vrgs_3$EN;

  // register vrgs_4
  reg [1 : 0] vrgs_4;
  wire [1 : 0] vrgs_4$D_IN;
  wire vrgs_4$EN;

  // register vrgs_5
  reg [1 : 0] vrgs_5;
  wire [1 : 0] vrgs_5$D_IN;
  wire vrgs_5$EN;

  // register vrgs_6
  reg [1 : 0] vrgs_6;
  wire [1 : 0] vrgs_6$D_IN;
  wire vrgs_6$EN;

  // register vrgs_7
  reg [1 : 0] vrgs_7;
  wire [1 : 0] vrgs_7$D_IN;
  wire vrgs_7$EN;

  // ports of submodule axis_xactor_f_data
  wire [760 : 0] axis_xactor_f_data$D_IN, axis_xactor_f_data$D_OUT;
  wire axis_xactor_f_data$CLR,
       axis_xactor_f_data$DEQ,
       axis_xactor_f_data$EMPTY_N,
       axis_xactor_f_data$ENQ,
       axis_xactor_f_data$FULL_N;

  // ports of submodule beatFF
  wire [31 : 0] beatFF$D_IN, beatFF$D_OUT;
  wire beatFF$CLR, beatFF$DEQ, beatFF$EMPTY_N, beatFF$ENQ, beatFF$FULL_N;

  // ports of submodule bridge_fIncomingData
  wire [31 : 0] bridge_fIncomingData$D_IN, bridge_fIncomingData$D_OUT;
  wire bridge_fIncomingData$CLR,
       bridge_fIncomingData$DEQ,
       bridge_fIncomingData$EMPTY_N,
       bridge_fIncomingData$ENQ,
       bridge_fIncomingData$FULL_N;

  // ports of submodule bridge_fOutgoingData
  wire [31 : 0] bridge_fOutgoingData$D_IN;
  wire bridge_fOutgoingData$CLR,
       bridge_fOutgoingData$DEQ,
       bridge_fOutgoingData$EMPTY_N,
       bridge_fOutgoingData$ENQ,
       bridge_fOutgoingData$FULL_N;

  // ports of submodule fOut_f
  wire [31 : 0] fOut_f$D_IN, fOut_f$D_OUT;
  wire fOut_f$CLR, fOut_f$DEQ, fOut_f$EMPTY_N, fOut_f$ENQ, fOut_f$FULL_N;

  // rule scheduling signals
  wire WILL_FIRE_RL_bridge_recv_beat_from_tcp,
       WILL_FIRE_RL_initializeBridge,
       WILL_FIRE_RL_xferBeat;

  // inputs to muxes for submodule ports
  wire [31 : 0] MUX_bridge_rFileHandle$write_1__VAL_1;

  // declarations used by system tasks
  // synopsys translate_off
  reg [135 : 0] TASK_bluenoc_recv_tcp_beat___d14;
  reg [7 : 0] b__h1134;
  reg [63 : 0] v__h1235;
  reg [31 : 0] b__h1366;
  // synopsys translate_on

  // remaining internal signals
  reg [31 : 0] x__h12556;
  wire [31 : 0] axis_xactor_f_dataD_OUT_BITS_760_TO_729_PLUS__ETC__q1,
		x__h11700;
  wire [7 : 0] IF_bridge_rBytesToTCP_0_EQ_0_1_THEN_4_ELSE_bri_ETC___d32,
	       bridge_rBytesFromTCP_PLUS_TASK_bluenoc_recv_tc_ETC___d16;
  wire cnt_1_EQ_vecSize_2___d63;

  // value method axi_in_m_tready
  assign axi_in_tready = axis_xactor_f_data$FULL_N || !tracesOn ;

  // submodule aresetAsserted
  ResetToBool aresetAsserted(.RST(RST_N_aresetn), .VAL());

  // submodule axis_xactor_f_data
  FIFO2 #(.width(32'd761),
	  .guarded(32'd1)) axis_xactor_f_data(.RST(RST_N_aresetn),
					      .CLK(CLK_aclk),
					      .D_IN(axis_xactor_f_data$D_IN),
					      .ENQ(axis_xactor_f_data$ENQ),
					      .DEQ(axis_xactor_f_data$DEQ),
					      .CLR(axis_xactor_f_data$CLR),
					      .D_OUT(axis_xactor_f_data$D_OUT),
					      .FULL_N(axis_xactor_f_data$FULL_N),
					      .EMPTY_N(axis_xactor_f_data$EMPTY_N));

  // submodule beatFF
  FIFO2 #(.width(32'd32), .guarded(32'd1)) beatFF(.RST(RST_N_aresetn),
						  .CLK(CLK_aclk),
						  .D_IN(beatFF$D_IN),
						  .ENQ(beatFF$ENQ),
						  .DEQ(beatFF$DEQ),
						  .CLR(beatFF$CLR),
						  .D_OUT(beatFF$D_OUT),
						  .FULL_N(beatFF$FULL_N),
						  .EMPTY_N(beatFF$EMPTY_N));

  // submodule bridge_fIncomingData
  FIFOL1 #(.width(32'd32)) bridge_fIncomingData(.RST(RST_N_aresetn),
						.CLK(CLK_aclk),
						.D_IN(bridge_fIncomingData$D_IN),
						.ENQ(bridge_fIncomingData$ENQ),
						.DEQ(bridge_fIncomingData$DEQ),
						.CLR(bridge_fIncomingData$CLR),
						.D_OUT(bridge_fIncomingData$D_OUT),
						.FULL_N(bridge_fIncomingData$FULL_N),
						.EMPTY_N(bridge_fIncomingData$EMPTY_N));

  // submodule bridge_fOutgoingData
  FIFOL1 #(.width(32'd32)) bridge_fOutgoingData(.RST(RST_N_aresetn),
						.CLK(CLK_aclk),
						.D_IN(bridge_fOutgoingData$D_IN),
						.ENQ(bridge_fOutgoingData$ENQ),
						.DEQ(bridge_fOutgoingData$DEQ),
						.CLR(bridge_fOutgoingData$CLR),
						.D_OUT(),
						.FULL_N(bridge_fOutgoingData$FULL_N),
						.EMPTY_N(bridge_fOutgoingData$EMPTY_N));

  // submodule fOut_f
  FIFO2 #(.width(32'd32), .guarded(32'd0)) fOut_f(.RST(RST_N_aresetn),
						  .CLK(CLK_aclk),
						  .D_IN(fOut_f$D_IN),
						  .ENQ(fOut_f$ENQ),
						  .DEQ(fOut_f$DEQ),
						  .CLR(fOut_f$CLR),
						  .D_OUT(fOut_f$D_OUT),
						  .FULL_N(fOut_f$FULL_N),
						  .EMPTY_N(fOut_f$EMPTY_N));

  // rule RL_xferBeat
  assign WILL_FIRE_RL_xferBeat =
	     beatFF$FULL_N &&
	     (!cnt_1_EQ_vecSize_2___d63 || axis_xactor_f_data$EMPTY_N) ;

  // rule RL_bridge_recv_beat_from_tcp
  assign WILL_FIRE_RL_bridge_recv_beat_from_tcp =
	     bridge_fOutgoingData$FULL_N && !bridge_rFileHandle[31] &&
	     (bridge_rBytesFromTCP == 8'd0 || bridge_rBytesFromTCP == 8'd4) ;

  // rule RL_initializeBridge
  assign WILL_FIRE_RL_initializeBridge =
	     bridge_rFileHandle == 32'hFFFFFFFF && !bridge_inReset_isInReset ;

  // inputs to muxes for submodule ports
  assign MUX_bridge_rFileHandle$write_1__VAL_1 =
	     b__h1366[31] ? 32'hFFFFFFFF : b__h1366 ;

  // inlined wires
  assign fOut_dst_ok$wget =
	     bridge_fIncomingData$FULL_N && !bridge_rFileHandle[31] ;

  // register bridge_inReset_isInReset
  assign bridge_inReset_isInReset$D_IN = 1'd0 ;
  assign bridge_inReset_isInReset$EN = bridge_inReset_isInReset ;

  // register bridge_rBeatFromTCP
  assign bridge_rBeatFromTCP$D_IN = TASK_bluenoc_recv_tcp_beat___d14[39:8] ;
  assign bridge_rBeatFromTCP$EN =
	     WILL_FIRE_RL_bridge_recv_beat_from_tcp &&
	     bridge_rBytesFromTCP_PLUS_TASK_bluenoc_recv_tc_ETC___d16 !=
	     8'd4 ;

  // register bridge_rBeatToTCP
  assign bridge_rBeatToTCP$D_IN = 32'h0 ;
  assign bridge_rBeatToTCP$EN = 1'b0 ;

  // register bridge_rBytesFromTCP
  assign bridge_rBytesFromTCP$D_IN =
	     (bridge_rBytesFromTCP_PLUS_TASK_bluenoc_recv_tc_ETC___d16 ==
	      8'd4) ?
	       8'd0 :
	       bridge_rBytesFromTCP_PLUS_TASK_bluenoc_recv_tc_ETC___d16 ;
  assign bridge_rBytesFromTCP$EN = WILL_FIRE_RL_bridge_recv_beat_from_tcp ;

  // register bridge_rBytesToTCP
  assign bridge_rBytesToTCP$D_IN =
	     (b__h1134 == 8'd4) ? 8'd0 : 8'd4 - b__h1134 ;
  assign bridge_rBytesToTCP$EN = bridge_fIncomingData$EMPTY_N ;

  // register bridge_rFileHandle
  assign bridge_rFileHandle$D_IN = MUX_bridge_rFileHandle$write_1__VAL_1 ;
  assign bridge_rFileHandle$EN = WILL_FIRE_RL_initializeBridge ;

  // register cnt
  assign cnt$D_IN = cnt_1_EQ_vecSize_2___d63 ? 8'd0 : cnt + 8'd1 ;
  assign cnt$EN = WILL_FIRE_RL_xferBeat ;

  // register trace
  assign trace$D_IN = axis_xactor_f_data$D_OUT[728:153] ;
  assign trace$EN = WILL_FIRE_RL_xferBeat && cnt_1_EQ_vecSize_2___d63 ;

  // register tracesOn
  assign tracesOn$D_IN = vrgs_0 == 2'd1 ;
  assign tracesOn$EN = vrgs_0 == 2'd1 || vrgs_0 == 2'd2 ;

  // register vecSize
  assign vecSize$D_IN =
	     axis_xactor_f_dataD_OUT_BITS_760_TO_729_PLUS__ETC__q1[7:0] ;
  assign vecSize$EN = WILL_FIRE_RL_xferBeat && cnt_1_EQ_vecSize_2___d63 ;

  // register vrgs_0
  assign vrgs_0$D_IN = vrgs_1 ;
  assign vrgs_0$EN = 1'd1 ;

  // register vrgs_1
  assign vrgs_1$D_IN = vrgs_2 ;
  assign vrgs_1$EN = 1'd1 ;

  // register vrgs_2
  assign vrgs_2$D_IN = vrgs_3 ;
  assign vrgs_2$EN = 1'd1 ;

  // register vrgs_3
  assign vrgs_3$D_IN = vrgs_4 ;
  assign vrgs_3$EN = 1'd1 ;

  // register vrgs_4
  assign vrgs_4$D_IN = vrgs_5 ;
  assign vrgs_4$EN = 1'd1 ;

  // register vrgs_5
  assign vrgs_5$D_IN = vrgs_6 ;
  assign vrgs_5$EN = 1'd1 ;

  // register vrgs_6
  assign vrgs_6$D_IN = vrgs_7 ;
  assign vrgs_6$EN = 1'd1 ;

  // register vrgs_7
  assign vrgs_7$D_IN = tvswitch ;
  assign vrgs_7$EN = 1'd1 ;

  // submodule axis_xactor_f_data
  assign axis_xactor_f_data$D_IN =
	     { axi_in_tdata, axi_in_tstrb, axi_in_tkeep, axi_in_tlast } ;
  assign axis_xactor_f_data$ENQ =
	     axi_in_tvalid && tracesOn && axis_xactor_f_data$FULL_N ;
  assign axis_xactor_f_data$DEQ =
	     WILL_FIRE_RL_xferBeat && cnt_1_EQ_vecSize_2___d63 ;
  assign axis_xactor_f_data$CLR = 1'b0 ;

  // submodule beatFF
  assign beatFF$D_IN = cnt_1_EQ_vecSize_2___d63 ? x__h11700 : x__h12556 ;
  assign beatFF$ENQ = WILL_FIRE_RL_xferBeat ;
  assign beatFF$DEQ = beatFF$EMPTY_N && fOut_f$FULL_N ;
  assign beatFF$CLR = 1'b0 ;

  // submodule bridge_fIncomingData
  assign bridge_fIncomingData$D_IN = fOut_f$D_OUT ;
  assign bridge_fIncomingData$ENQ =
	     bridge_fIncomingData$FULL_N && fOut_f$EMPTY_N ;
  assign bridge_fIncomingData$DEQ =
	     bridge_fIncomingData$EMPTY_N && b__h1134 == 8'd4 ;
  assign bridge_fIncomingData$CLR = 1'b0 ;

  // submodule bridge_fOutgoingData
  assign bridge_fOutgoingData$D_IN = TASK_bluenoc_recv_tcp_beat___d14[39:8] ;
  assign bridge_fOutgoingData$ENQ =
	     WILL_FIRE_RL_bridge_recv_beat_from_tcp &&
	     bridge_rBytesFromTCP_PLUS_TASK_bluenoc_recv_tc_ETC___d16 ==
	     8'd4 ;
  assign bridge_fOutgoingData$DEQ = bridge_fOutgoingData$EMPTY_N ;
  assign bridge_fOutgoingData$CLR = 1'b0 ;

  // submodule fOut_f
  assign fOut_f$D_IN = beatFF$D_OUT ;
  assign fOut_f$ENQ = beatFF$EMPTY_N && fOut_f$FULL_N ;
  assign fOut_f$DEQ = fOut_f$EMPTY_N && fOut_dst_ok$wget ;
  assign fOut_f$CLR = 1'b0 ;

  // remaining internal signals
  assign IF_bridge_rBytesToTCP_0_EQ_0_1_THEN_4_ELSE_bri_ETC___d32 =
	     (bridge_rBytesToTCP == 8'd0) ? 8'd4 : bridge_rBytesToTCP ;
  assign axis_xactor_f_dataD_OUT_BITS_760_TO_729_PLUS__ETC__q1 =
	     (axis_xactor_f_data$D_OUT[760:729] + 32'd4 - 32'd1) >> 2 ;
  assign bridge_rBytesFromTCP_PLUS_TASK_bluenoc_recv_tc_ETC___d16 =
	     bridge_rBytesFromTCP + TASK_bluenoc_recv_tcp_beat___d14[7:0] ;
  assign cnt_1_EQ_vecSize_2___d63 = cnt == vecSize ;
  assign x__h11700 = { 8'd1, axis_xactor_f_data$D_OUT[736:729], 16'd256 } ;
  always@(cnt or trace)
  begin
    case (cnt)
      8'd0: x__h12556 = trace[31:0];
      8'd1: x__h12556 = trace[63:32];
      8'd2: x__h12556 = trace[95:64];
      8'd3: x__h12556 = trace[127:96];
      8'd4: x__h12556 = trace[159:128];
      8'd5: x__h12556 = trace[191:160];
      8'd6: x__h12556 = trace[223:192];
      8'd7: x__h12556 = trace[255:224];
      8'd8: x__h12556 = trace[287:256];
      8'd9: x__h12556 = trace[319:288];
      8'd10: x__h12556 = trace[351:320];
      8'd11: x__h12556 = trace[383:352];
      8'd12: x__h12556 = trace[415:384];
      8'd13: x__h12556 = trace[447:416];
      8'd14: x__h12556 = trace[479:448];
      8'd15: x__h12556 = trace[511:480];
      8'd16: x__h12556 = trace[543:512];
      8'd17: x__h12556 = trace[575:544];
      default: x__h12556 = 32'hAAAAAAAA /* unspecified value */ ;
    endcase
  end

  // handling of inlined registers

  always@(posedge CLK_aclk)
  begin
    if (RST_N_aresetn == `BSV_RESET_VALUE)
      begin
        bridge_rBytesFromTCP <= `BSV_ASSIGNMENT_DELAY 8'd0;
	bridge_rBytesToTCP <= `BSV_ASSIGNMENT_DELAY 8'd0;
	bridge_rFileHandle <= `BSV_ASSIGNMENT_DELAY 32'hFFFFFFFF;
	cnt <= `BSV_ASSIGNMENT_DELAY 8'd0;
	tracesOn <= `BSV_ASSIGNMENT_DELAY 1'd0;
	vecSize <= `BSV_ASSIGNMENT_DELAY 8'd0;
	vrgs_0 <= `BSV_ASSIGNMENT_DELAY 2'd0;
	vrgs_1 <= `BSV_ASSIGNMENT_DELAY 2'd0;
	vrgs_2 <= `BSV_ASSIGNMENT_DELAY 2'd0;
	vrgs_3 <= `BSV_ASSIGNMENT_DELAY 2'd0;
	vrgs_4 <= `BSV_ASSIGNMENT_DELAY 2'd0;
	vrgs_5 <= `BSV_ASSIGNMENT_DELAY 2'd0;
	vrgs_6 <= `BSV_ASSIGNMENT_DELAY 2'd0;
	vrgs_7 <= `BSV_ASSIGNMENT_DELAY 2'd0;
      end
    else
      begin
        if (bridge_rBytesFromTCP$EN)
	  bridge_rBytesFromTCP <= `BSV_ASSIGNMENT_DELAY
	      bridge_rBytesFromTCP$D_IN;
	if (bridge_rBytesToTCP$EN)
	  bridge_rBytesToTCP <= `BSV_ASSIGNMENT_DELAY bridge_rBytesToTCP$D_IN;
	if (bridge_rFileHandle$EN)
	  bridge_rFileHandle <= `BSV_ASSIGNMENT_DELAY bridge_rFileHandle$D_IN;
	if (cnt$EN) cnt <= `BSV_ASSIGNMENT_DELAY cnt$D_IN;
	if (tracesOn$EN) tracesOn <= `BSV_ASSIGNMENT_DELAY tracesOn$D_IN;
	if (vecSize$EN) vecSize <= `BSV_ASSIGNMENT_DELAY vecSize$D_IN;
	if (vrgs_0$EN) vrgs_0 <= `BSV_ASSIGNMENT_DELAY vrgs_0$D_IN;
	if (vrgs_1$EN) vrgs_1 <= `BSV_ASSIGNMENT_DELAY vrgs_1$D_IN;
	if (vrgs_2$EN) vrgs_2 <= `BSV_ASSIGNMENT_DELAY vrgs_2$D_IN;
	if (vrgs_3$EN) vrgs_3 <= `BSV_ASSIGNMENT_DELAY vrgs_3$D_IN;
	if (vrgs_4$EN) vrgs_4 <= `BSV_ASSIGNMENT_DELAY vrgs_4$D_IN;
	if (vrgs_5$EN) vrgs_5 <= `BSV_ASSIGNMENT_DELAY vrgs_5$D_IN;
	if (vrgs_6$EN) vrgs_6 <= `BSV_ASSIGNMENT_DELAY vrgs_6$D_IN;
	if (vrgs_7$EN) vrgs_7 <= `BSV_ASSIGNMENT_DELAY vrgs_7$D_IN;
      end
    if (bridge_rBeatFromTCP$EN)
      bridge_rBeatFromTCP <= `BSV_ASSIGNMENT_DELAY bridge_rBeatFromTCP$D_IN;
    if (bridge_rBeatToTCP$EN)
      bridge_rBeatToTCP <= `BSV_ASSIGNMENT_DELAY bridge_rBeatToTCP$D_IN;
    if (trace$EN) trace <= `BSV_ASSIGNMENT_DELAY trace$D_IN;
  end

  always@(posedge CLK_aclk or `BSV_RESET_EDGE RST_N_aresetn)
  if (RST_N_aresetn == `BSV_RESET_VALUE)
    begin
      bridge_inReset_isInReset <= `BSV_ASSIGNMENT_DELAY 1'd1;
    end
  else
    begin
      if (bridge_inReset_isInReset$EN)
	bridge_inReset_isInReset <= `BSV_ASSIGNMENT_DELAY
	    bridge_inReset_isInReset$D_IN;
    end

  // synopsys translate_off
  `ifdef BSV_NO_INITIAL_BLOCKS
  `else // not BSV_NO_INITIAL_BLOCKS
  initial
  begin
    bridge_inReset_isInReset = 1'h0;
    bridge_rBeatFromTCP = 32'hAAAAAAAA;
    bridge_rBeatToTCP = 32'hAAAAAAAA;
    bridge_rBytesFromTCP = 8'hAA;
    bridge_rBytesToTCP = 8'hAA;
    bridge_rFileHandle = 32'hAAAAAAAA;
    cnt = 8'hAA;
    trace =
	576'hAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA;
    tracesOn = 1'h0;
    vecSize = 8'hAA;
    vrgs_0 = 2'h2;
    vrgs_1 = 2'h2;
    vrgs_2 = 2'h2;
    vrgs_3 = 2'h2;
    vrgs_4 = 2'h2;
    vrgs_5 = 2'h2;
    vrgs_6 = 2'h2;
    vrgs_7 = 2'h2;
  end
  `endif // BSV_NO_INITIAL_BLOCKS
  // synopsys translate_on

  // handling of system tasks

  // synopsys translate_off
  always@(negedge CLK_aclk)
  begin
    #0;
    if (RST_N_aresetn != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_bridge_recv_beat_from_tcp)
	begin
	   bluenoc_recv_tcp_beat(TASK_bluenoc_recv_tcp_beat___d14,
				 bridge_rFileHandle,
				 8'd4,
				 bridge_rBytesFromTCP,
				 { 96'd0, bridge_rBeatFromTCP });
	  #0;
	end
    if (RST_N_aresetn != `BSV_RESET_VALUE)
      if (bridge_fIncomingData$EMPTY_N)
	begin
	  b__h1134 =
	      bluenoc_send_tcp_beat(bridge_rFileHandle,
					      8'd4,
					      IF_bridge_rBytesToTCP_0_EQ_0_1_THEN_4_ELSE_bri_ETC___d32,
					      { 96'd0,
						bridge_fIncomingData$D_OUT });
	  #0;
	end
    if (RST_N_aresetn != `BSV_RESET_VALUE)
      if (bridge_fIncomingData$EMPTY_N && b__h1134 == 8'd4)
	begin
	  v__h1235 = $time;
	  #0;
	end
    if (RST_N_aresetn != `BSV_RESET_VALUE)
      if (bridge_fIncomingData$EMPTY_N && b__h1134 == 8'd4)
	$display("[%t] HW_SEND %d %x",
		 v__h1235,
		 $unsigned(IF_bridge_rBytesToTCP_0_EQ_0_1_THEN_4_ELSE_bri_ETC___d32),
		 bridge_fIncomingData$D_OUT);
    if (RST_N_aresetn != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_initializeBridge)
	begin
	  b__h1366 = bluenoc_open_tcp_socket(32'h0000357B);
	  #0;
	end
    if (RST_N_aresetn != `BSV_RESET_VALUE)
      if (WILL_FIRE_RL_initializeBridge && b__h1366[31])
	$display("Couldn't listen!");
  end
  // synopsys translate_on
endmodule  // mkSVF_Bridge
